magic
tech sky130A
timestamp 1670170588
<< nmos >>
rect 0 -95 15 10
<< ndiff >>
rect -60 -95 0 10
rect 15 -95 75 10
<< poly >>
rect 0 10 15 25
rect 0 -110 15 -95
<< locali >>
rect -50 -85 -10 0
rect 25 -85 65 0
<< end >>
